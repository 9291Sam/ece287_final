module random(input clk, output reg[255:0] rand);

// python :)
always @ (posedge clk)
    rand <= 
        255'b0101111101001000111000110000011111111011011111111001111111001000011111110111111011001000111110010101110000111111000101110010110110100011010111010111111101010111000100100110100010010101101010001111011000111001111000111111001110101011101110110111110110100100
        + {
        rand[93] ^ /* ~ */ rand[81] ^ rand[143],
        rand[33] ^ /* ~ */ rand[73] ^ rand[243],
        rand[94] ^ /* ~ */ rand[165] ^ rand[125],
        rand[172] ^ /* ~ */ rand[220] ^ rand[23],
        rand[248] ^ /* ~ */ rand[79] ^ rand[177],
        rand[44] ^ /* ~ */ rand[216] ^ rand[185],
        rand[108] ^ /* ~ */ rand[130] ^ rand[15],
        rand[53] ^ /* ~ */ rand[164] ^ rand[9],
        rand[60] ^ /* ~ */ rand[101] ^ rand[13],
        rand[198] ^ /* ~ */ rand[1] ^ rand[13],
        rand[156] ^ /* ~ */ rand[208] ^ rand[94],
        rand[65] ^ /* ~ */ rand[160] ^ rand[85],
        rand[172] ^ /* ~ */ rand[152] ^ rand[197],
        rand[241] ^ /* ~ */ rand[45] ^ rand[146],
        rand[225] ^ /* ~ */ rand[175] ^ rand[33],
        rand[185] ^ /* ~ */ rand[144] ^ rand[241],
        rand[152] ^ /* ~ */ rand[96] ^ rand[155],
        rand[114] ^ /* ~ */ rand[99] ^ rand[97],
        rand[196] ^ /* ~ */ rand[228] ^ rand[13],
        rand[206] ^ /* ~ */ rand[198] ^ rand[180],
        rand[125] ^ /* ~ */ rand[209] ^ rand[40],
        rand[119] ^ /* ~ */ rand[82] ^ rand[35],
        rand[159] ^ /* ~ */ rand[101] ^ rand[174],
        rand[254] ^ /* ~ */ rand[23] ^ rand[247],
        rand[229] ^ /* ~ */ rand[78] ^ rand[12],
        rand[28] ^ /* ~ */ rand[58] ^ rand[63],
        rand[45] ^ /* ~ */ rand[126] ^ rand[213],
        rand[75] ^ /* ~ */ rand[183] ^ rand[56],
        rand[195] ^ /* ~ */ rand[118] ^ rand[199],
        rand[233] ^ /* ~ */ rand[129] ^ rand[29],
        rand[67] ^ /* ~ */ rand[28] ^ rand[215],
        rand[114] ^ /* ~ */ rand[81] ^ rand[89],
        rand[46] ^ /* ~ */ rand[60] ^ rand[196],
        rand[185] ^ /* ~ */ rand[35] ^ rand[126],
        rand[230] ^ /* ~ */ rand[147] ^ rand[168],
        rand[177] ^ /* ~ */ rand[111] ^ rand[61],
        rand[130] ^ /* ~ */ rand[241] ^ rand[123],
        rand[64] ^ /* ~ */ rand[65] ^ rand[42],
        rand[119] ^ /* ~ */ rand[35] ^ rand[29],
        rand[178] ^ /* ~ */ rand[42] ^ rand[7],
        rand[159] ^ /* ~ */ rand[79] ^ rand[79],
        rand[21] ^ /* ~ */ rand[201] ^ rand[57],
        rand[141] ^ /* ~ */ rand[189] ^ rand[63],
        rand[103] ^ /* ~ */ rand[216] ^ rand[32],
        rand[0] ^ /* ~ */ rand[7] ^ rand[157],
        rand[114] ^ /* ~ */ rand[8] ^ rand[188],
        rand[46] ^ /* ~ */ rand[194] ^ rand[197],
        rand[206] ^ /* ~ */ rand[47] ^ rand[225],
        rand[208] ^ /* ~ */ rand[200] ^ rand[156],
        rand[232] ^ /* ~ */ rand[252] ^ rand[132],
        rand[211] ^ /* ~ */ rand[68] ^ rand[214],
        rand[65] ^ /* ~ */ rand[195] ^ rand[183],
        rand[64] ^ /* ~ */ rand[213] ^ rand[139],
        rand[146] ^ /* ~ */ rand[116] ^ rand[234],
        rand[177] ^ /* ~ */ rand[187] ^ rand[66],
        rand[121] ^ /* ~ */ rand[252] ^ rand[136],
        rand[183] ^ /* ~ */ rand[206] ^ rand[19],
        rand[169] ^ /* ~ */ rand[181] ^ rand[236],
        rand[193] ^ /* ~ */ rand[231] ^ rand[157],
        rand[39] ^ /* ~ */ rand[89] ^ rand[176],
        rand[112] ^ /* ~ */ rand[18] ^ rand[184],
        rand[111] ^ /* ~ */ rand[133] ^ rand[52],
        rand[216] ^ /* ~ */ rand[126] ^ rand[251],
        rand[192] ^ /* ~ */ rand[145] ^ rand[82],
        rand[138] ^ /* ~ */ rand[57] ^ rand[196],
        rand[68] ^ /* ~ */ rand[59] ^ rand[236],
        rand[12] ^ /* ~ */ rand[12] ^ rand[17],
        rand[166] ^ /* ~ */ rand[162] ^ rand[56],
        rand[101] ^ /* ~ */ rand[127] ^ rand[140],
        rand[156] ^ /* ~ */ rand[61] ^ rand[91],
        rand[7] ^ /* ~ */ rand[202] ^ rand[68],
        rand[141] ^ /* ~ */ rand[111] ^ rand[59],
        rand[177] ^ /* ~ */ rand[26] ^ rand[192],
        rand[83] ^ /* ~ */ rand[10] ^ rand[141],
        rand[32] ^ /* ~ */ rand[235] ^ rand[152],
        rand[109] ^ /* ~ */ rand[222] ^ rand[205],
        rand[212] ^ /* ~ */ rand[39] ^ rand[78],
        rand[44] ^ /* ~ */ rand[239] ^ rand[249],
        rand[192] ^ /* ~ */ rand[155] ^ rand[51],
        rand[206] ^ /* ~ */ rand[13] ^ rand[251],
        rand[166] ^ /* ~ */ rand[0] ^ rand[192],
        rand[82] ^ /* ~ */ rand[70] ^ rand[21],
        rand[8] ^ /* ~ */ rand[31] ^ rand[148],
        rand[190] ^ /* ~ */ rand[136] ^ rand[114],
        rand[205] ^ /* ~ */ rand[73] ^ rand[252],
        rand[241] ^ /* ~ */ rand[96] ^ rand[173],
        rand[17] ^ /* ~ */ rand[83] ^ rand[185],
        rand[192] ^ /* ~ */ rand[47] ^ rand[113],
        rand[30] ^ /* ~ */ rand[12] ^ rand[201],
        rand[84] ^ /* ~ */ rand[216] ^ rand[252],
        rand[96] ^ /* ~ */ rand[235] ^ rand[66],
        rand[189] ^ /* ~ */ rand[139] ^ rand[95],
        rand[184] ^ /* ~ */ rand[8] ^ rand[209],
        rand[47] ^ /* ~ */ rand[195] ^ rand[10],
        rand[37] ^ /* ~ */ rand[8] ^ rand[53],
        rand[9] ^ /* ~ */ rand[186] ^ rand[81],
        rand[210] ^ /* ~ */ rand[1] ^ rand[42],
        rand[193] ^ /* ~ */ rand[215] ^ rand[83],
        rand[3] ^ /* ~ */ rand[74] ^ rand[243],
        rand[95] ^ /* ~ */ rand[119] ^ rand[80],
        rand[9] ^ /* ~ */ rand[163] ^ rand[160],
        rand[221] ^ /* ~ */ rand[98] ^ rand[127],
        rand[48] ^ /* ~ */ rand[236] ^ rand[244],
        rand[199] ^ /* ~ */ rand[144] ^ rand[128],
        rand[146] ^ /* ~ */ rand[12] ^ rand[184],
        rand[156] ^ /* ~ */ rand[126] ^ rand[232],
        rand[51] ^ /* ~ */ rand[92] ^ rand[220],
        rand[62] ^ /* ~ */ rand[198] ^ rand[126],
        rand[247] ^ /* ~ */ rand[250] ^ rand[17],
        rand[248] ^ /* ~ */ rand[102] ^ rand[244],
        rand[240] ^ /* ~ */ rand[145] ^ rand[109],
        rand[152] ^ /* ~ */ rand[56] ^ rand[250],
        rand[119] ^ /* ~ */ rand[1] ^ rand[146],
        rand[47] ^ /* ~ */ rand[72] ^ rand[249],
        rand[135] ^ /* ~ */ rand[170] ^ rand[22],
        rand[215] ^ /* ~ */ rand[159] ^ rand[107],
        rand[87] ^ /* ~ */ rand[172] ^ rand[174],
        rand[206] ^ /* ~ */ rand[120] ^ rand[228],
        rand[176] ^ /* ~ */ rand[230] ^ rand[224],
        rand[144] ^ /* ~ */ rand[206] ^ rand[11],
        rand[116] ^ /* ~ */ rand[93] ^ rand[191],
        rand[40] ^ /* ~ */ rand[37] ^ rand[133],
        rand[36] ^ /* ~ */ rand[236] ^ rand[192],
        rand[219] ^ /* ~ */ rand[111] ^ rand[58],
        rand[3] ^ /* ~ */ rand[175] ^ rand[235],
        rand[180] ^ /* ~ */ rand[7] ^ rand[115],
        rand[82] ^ /* ~ */ rand[96] ^ rand[167],
        rand[252] ^ /* ~ */ rand[4] ^ rand[89],
        rand[226] ^ /* ~ */ rand[51] ^ rand[117],
        rand[103] ^ /* ~ */ rand[146] ^ rand[121],
        rand[186] ^ /* ~ */ rand[44] ^ rand[5],
        rand[173] ^ /* ~ */ rand[231] ^ rand[64],
        rand[25] ^ /* ~ */ rand[165] ^ rand[37],
        rand[0] ^ /* ~ */ rand[24] ^ rand[130],
        rand[80] ^ /* ~ */ rand[126] ^ rand[68],
        rand[112] ^ /* ~ */ rand[86] ^ rand[32],
        rand[107] ^ /* ~ */ rand[140] ^ rand[50],
        rand[138] ^ /* ~ */ rand[112] ^ rand[132],
        rand[54] ^ /* ~ */ rand[78] ^ rand[69],
        rand[177] ^ /* ~ */ rand[109] ^ rand[136],
        rand[206] ^ /* ~ */ rand[234] ^ rand[214],
        rand[232] ^ /* ~ */ rand[252] ^ rand[77],
        rand[153] ^ /* ~ */ rand[78] ^ rand[62],
        rand[85] ^ /* ~ */ rand[157] ^ rand[17],
        rand[189] ^ /* ~ */ rand[252] ^ rand[14],
        rand[230] ^ /* ~ */ rand[41] ^ rand[157],
        rand[16] ^ /* ~ */ rand[186] ^ rand[4],
        rand[10] ^ /* ~ */ rand[198] ^ rand[205],
        rand[149] ^ /* ~ */ rand[125] ^ rand[0],
        rand[185] ^ /* ~ */ rand[141] ^ rand[129],
        rand[192] ^ /* ~ */ rand[82] ^ rand[27],
        rand[153] ^ /* ~ */ rand[144] ^ rand[237],
        rand[149] ^ /* ~ */ rand[207] ^ rand[190],
        rand[121] ^ /* ~ */ rand[195] ^ rand[244],
        rand[111] ^ /* ~ */ rand[69] ^ rand[61],
        rand[205] ^ /* ~ */ rand[206] ^ rand[130],
        rand[19] ^ /* ~ */ rand[239] ^ rand[39],
        rand[38] ^ /* ~ */ rand[205] ^ rand[208],
        rand[113] ^ /* ~ */ rand[60] ^ rand[32],
        rand[74] ^ /* ~ */ rand[254] ^ rand[85],
        rand[54] ^ /* ~ */ rand[150] ^ rand[133],
        rand[234] ^ /* ~ */ rand[5] ^ rand[70],
        rand[115] ^ /* ~ */ rand[220] ^ rand[191],
        rand[5] ^ /* ~ */ rand[204] ^ rand[196],
        rand[119] ^ /* ~ */ rand[200] ^ rand[223],
        rand[236] ^ /* ~ */ rand[123] ^ rand[211],
        rand[170] ^ /* ~ */ rand[59] ^ rand[170],
        rand[74] ^ /* ~ */ rand[156] ^ rand[166],
        rand[160] ^ /* ~ */ rand[130] ^ rand[182],
        rand[195] ^ /* ~ */ rand[236] ^ rand[36],
        rand[158] ^ /* ~ */ rand[21] ^ rand[158],
        rand[91] ^ /* ~ */ rand[91] ^ rand[34],
        rand[117] ^ /* ~ */ rand[238] ^ rand[21],
        rand[244] ^ /* ~ */ rand[110] ^ rand[176],
        rand[125] ^ /* ~ */ rand[3] ^ rand[22],
        rand[70] ^ /* ~ */ rand[189] ^ rand[209],
        rand[72] ^ /* ~ */ rand[97] ^ rand[228],
        rand[67] ^ /* ~ */ rand[197] ^ rand[15],
        rand[24] ^ /* ~ */ rand[149] ^ rand[244],
        rand[13] ^ /* ~ */ rand[203] ^ rand[126],
        rand[253] ^ /* ~ */ rand[200] ^ rand[220],
        rand[131] ^ /* ~ */ rand[146] ^ rand[90],
        rand[74] ^ /* ~ */ rand[214] ^ rand[73],
        rand[28] ^ /* ~ */ rand[111] ^ rand[205],
        rand[199] ^ /* ~ */ rand[76] ^ rand[148],
        rand[90] ^ /* ~ */ rand[131] ^ rand[104],
        rand[11] ^ /* ~ */ rand[207] ^ rand[67],
        rand[27] ^ /* ~ */ rand[17] ^ rand[204],
        rand[60] ^ /* ~ */ rand[8] ^ rand[245],
        rand[238] ^ /* ~ */ rand[138] ^ rand[28],
        rand[104] ^ /* ~ */ rand[108] ^ rand[221],
        rand[119] ^ /* ~ */ rand[173] ^ rand[96],
        rand[2] ^ /* ~ */ rand[139] ^ rand[196],
        rand[6] ^ /* ~ */ rand[167] ^ rand[59],
        rand[126] ^ /* ~ */ rand[29] ^ rand[67],
        rand[218] ^ /* ~ */ rand[123] ^ rand[0],
        rand[123] ^ /* ~ */ rand[115] ^ rand[27],
        rand[36] ^ /* ~ */ rand[186] ^ rand[80],
        rand[212] ^ /* ~ */ rand[109] ^ rand[201],
        rand[101] ^ /* ~ */ rand[154] ^ rand[146],
        rand[200] ^ /* ~ */ rand[111] ^ rand[239],
        rand[57] ^ /* ~ */ rand[134] ^ rand[230],
        rand[63] ^ /* ~ */ rand[175] ^ rand[193],
        rand[88] ^ /* ~ */ rand[30] ^ rand[2],
        rand[81] ^ /* ~ */ rand[254] ^ rand[241],
        rand[92] ^ /* ~ */ rand[129] ^ rand[14],
        rand[107] ^ /* ~ */ rand[237] ^ rand[43],
        rand[73] ^ /* ~ */ rand[34] ^ rand[223],
        rand[143] ^ /* ~ */ rand[146] ^ rand[96],
        rand[135] ^ /* ~ */ rand[244] ^ rand[68],
        rand[211] ^ /* ~ */ rand[99] ^ rand[32],
        rand[61] ^ /* ~ */ rand[108] ^ rand[145],
        rand[194] ^ /* ~ */ rand[153] ^ rand[108],
        rand[197] ^ /* ~ */ rand[203] ^ rand[244],
        rand[106] ^ /* ~ */ rand[116] ^ rand[64],
        rand[114] ^ /* ~ */ rand[189] ^ rand[56],
        rand[242] ^ /* ~ */ rand[215] ^ rand[186],
        rand[21] ^ /* ~ */ rand[22] ^ rand[65],
        rand[251] ^ /* ~ */ rand[234] ^ rand[226],
        rand[243] ^ /* ~ */ rand[132] ^ rand[91],
        rand[29] ^ /* ~ */ rand[46] ^ rand[153],
        rand[24] ^ /* ~ */ rand[14] ^ rand[241],
        rand[148] ^ /* ~ */ rand[227] ^ rand[198],
        rand[149] ^ /* ~ */ rand[198] ^ rand[139],
        rand[134] ^ /* ~ */ rand[89] ^ rand[27],
        rand[193] ^ /* ~ */ rand[187] ^ rand[56],
        rand[51] ^ /* ~ */ rand[1] ^ rand[169],
        rand[250] ^ /* ~ */ rand[35] ^ rand[81],
        rand[41] ^ /* ~ */ rand[208] ^ rand[165],
        rand[193] ^ /* ~ */ rand[35] ^ rand[145],
        rand[151] ^ /* ~ */ rand[29] ^ rand[28],
        rand[30] ^ /* ~ */ rand[243] ^ rand[16],
        rand[180] ^ /* ~ */ rand[120] ^ rand[147],
        rand[136] ^ /* ~ */ rand[81] ^ rand[70],
        rand[192] ^ /* ~ */ rand[14] ^ rand[10],
        rand[224] ^ /* ~ */ rand[203] ^ rand[103],
        rand[247] ^ /* ~ */ rand[228] ^ rand[68],
        rand[50] ^ /* ~ */ rand[77] ^ rand[155],
        rand[49] ^ /* ~ */ rand[113] ^ rand[24],
        rand[139] ^ /* ~ */ rand[91] ^ rand[153],
        rand[5] ^ /* ~ */ rand[246] ^ rand[6],
        rand[38] ^ /* ~ */ rand[37] ^ rand[48],
        rand[34] ^ /* ~ */ rand[193] ^ rand[214],
        rand[53] ^ /* ~ */ rand[126] ^ rand[12],
        rand[175] ^ /* ~ */ rand[5] ^ rand[191],
        rand[94] ^ /* ~ */ rand[166] ^ rand[62],
        rand[167] ^ /* ~ */ rand[110] ^ rand[8],
        rand[221] ^ /* ~ */ rand[189] ^ rand[46],
        rand[148] ^ /* ~ */ rand[201] ^ rand[41],
        rand[53] ^ /* ~ */ rand[237] ^ rand[187],
        rand[72] ^ /* ~ */ rand[208] ^ rand[202],
        rand[187] ^ /* ~ */ rand[167] ^ rand[60],
        rand[134] ^ /* ~ */ rand[121] ^ rand[30],
        rand[162] ^ /* ~ */ rand[104] ^ rand[237],
        rand[170] ^ /* ~ */ rand[44] ^ rand[84]
    };


endmodule